* /home/nithish/Desktop/eSim/Examples/High_Pass_Filter/High_Pass_Filter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 14 Jun 2023 05:25:44 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  out GND 1k		
C1  out in 10u		
v1  in GND AC		
U1  in plot_v1		
U3  out plot_v1		

.end
