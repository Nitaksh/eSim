* /home/nithish/Desktop/eSim/Examples/Astable555/Astable555.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue 13 Jun 2023 02:53:16 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R3  V_Out GND 1k		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 1k		
R2  Net-_R1-Pad2_ C_Out 10k		
v1  Net-_R1-Pad1_ GND DC		
C1  C_Out GND 0.1u		
C2  Net-_C2-Pad1_ GND 0.01u		
U2  V_Out plot_v1		
U1  C_Out plot_v1		
X1  GND C_Out V_Out Net-_R1-Pad1_ Net-_C2-Pad1_ C_Out Net-_R1-Pad2_ Net-_R1-Pad1_ LM555N		

.end
